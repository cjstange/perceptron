`default_nettype none 